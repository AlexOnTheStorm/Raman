library verilog;
use verilog.vl_types.all;
entity Raman is
    port(
        enable          : in     vl_logic;
        clk             : in     vl_logic;
        data            : in     vl_logic_vector(11 downto 0);
        ready           : out    vl_logic;
        ratio_enable    : out    vl_logic;
        start           : out    vl_logic;
        C0              : out    vl_logic;
        wrreq           : out    vl_logic;
        rdreq           : out    vl_logic;
        switch          : out    vl_logic;
        div_enable      : out    vl_logic;
        wren            : out    vl_logic;
        aclr            : out    vl_logic;
        wren_stokes     : out    vl_logic;
        wren_antistokes : out    vl_logic;
        wren_storage    : out    vl_logic;
        wren_temp       : out    vl_logic;
        cnt_div         : out    vl_logic_vector(10 downto 0);
        cnt_measure     : out    vl_logic_vector(16 downto 0);
        cnt_point       : out    vl_logic_vector(10 downto 0);
        cnt_ratio       : out    vl_logic_vector(10 downto 0);
        cnt_save        : out    vl_logic_vector(3 downto 0);
        datamem         : out    vl_logic_vector(28 downto 0);
        q               : out    vl_logic_vector(11 downto 0);
        q_storage       : out    vl_logic_vector(11 downto 0);
        qantistokes     : out    vl_logic_vector(28 downto 0);
        qout            : out    vl_logic_vector(11 downto 0);
        qstokes         : out    vl_logic_vector(28 downto 0);
        qsummary        : out    vl_logic_vector(28 downto 0);
        quot_ratio      : out    vl_logic_vector(11 downto 0);
        quotient        : out    vl_logic_vector(11 downto 0);
        rd_address_storage: out    vl_logic_vector(14 downto 0);
        rdaddress       : out    vl_logic_vector(10 downto 0);
        wr_address_storage: out    vl_logic_vector(14 downto 0);
        wraddr          : out    vl_logic_vector(10 downto 0)
    );
end Raman;
