library verilog;
use verilog.vl_types.all;
entity tbRam is
end tbRam;
