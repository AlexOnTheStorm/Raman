library verilog;
use verilog.vl_types.all;
entity MEASURES is
    port(
        result          : out    vl_logic_vector(16 downto 0)
    );
end MEASURES;
