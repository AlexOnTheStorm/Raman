library verilog;
use verilog.vl_types.all;
entity POINTS is
    port(
        result          : out    vl_logic_vector(10 downto 0)
    );
end POINTS;
